/*

*/
module top
(
    input CLK_12MHZ
);



endmodule